module AES_Encrypt(
	

)
